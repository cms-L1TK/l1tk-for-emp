library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.BDTTypes.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((5, 2, 5, 5, 4, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 5, 5, 4, 4, 6, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 2, 4, 4, 6, 6, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 6, 5, 4, 0, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 2, 4, 6, 4, 6, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 4, 5, 6, 5, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 4, 6, 6, 5, 5, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 4, 3, 6, 2, 2, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 4, 4, 6, 4, 6, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 4, 0, 6, 3, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 5, 5, 2, 2, -2, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 5, 5, 0, -2, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 4, 5, 0, 6, -2, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 4, 6, 6, 1, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 6, 5, 4, 2, 6, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 1, 5, 4, 0, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 5, 1, 0, -2, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 1, 1, 0, 0, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 5, 1, 4, 0, 0, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 1, 0, 1, 6, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 5, 0, 0, -2, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 0, 0, 5, 0, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 5, 2, 1, 1, 1, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 0, 0, 1, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 0, 1, 0, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 4, 5, 0, 1, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 1, 1, 1, 0, -2, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 0, 6, 6, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 6, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 5, -2, 6, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 0, 5, 0, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 0, 6, 1, 0, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 1, 0, -2, 1, 5, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 6, 0, 1, 2, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 1, 1, 2, 5, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 1, 0, 1, 1, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 4, 6, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 6, 0, 4, 6, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 0, 1, 4, 0, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 0, -2, 6, 6, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 0, 1, -2, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 1, 0, 4, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 6, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 0, 0, 0, 0, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 1, 1, 1, 1, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 6, 6, 1, 1, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 5, 1, 0, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 2, 1, 0, -2, 5, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 5, 0, 1, 2, 5, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 0, 1, 1, -2, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 6, 1, 4, 6, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 4, 0, 6, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 1, 1, 0, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 0, 1, 2, 0, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 4, 6, 5, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 0, 0, 0, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 6, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 5, 4, -2, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 1, 1, 2, 1, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 0, 1, 1, -2, 0, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((304, 144, 400, 272, 48, 48, 16, 0, 0, 0, 0, 0, 0, 0, 0),
                (336, 272, 464, 48, 48, 304, -54, 0, 0, 0, 0, 0, 0, 0, 0),
                (304, 144, 16, 48, 112, 272, 432, 0, 0, 0, 0, 0, 0, 0, 0),
                (272, 368, 432, 48, 32, 112, 144, 0, 0, 0, 0, 0, 0, 0, 0),
                (272, 144, 16, 368, 16, 144, 112, 0, 0, 0, 0, 0, 0, 0, 0),
                (336, 16, 464, 304, 112, 48, -54, 0, 0, 0, 0, 0, 0, 0, 0),
                (240, 48, 432, 304, 48, 464, 16, 0, 0, 0, 0, 0, 0, 0, 0),
                (208, 16, 144, 304, 112, 144, 208, 0, 0, 0, 0, 0, 0, 0, 0),
                (176, 48, 16, 304, 80, 208, 80, 0, 0, 0, 0, 0, 0, 0, 0),
                (336, 16, 57, 208, 144, -56, -11, 0, 0, 0, 0, 0, 0, 0, 0),
                (144, 112, 432, 80, 48, 0, 48, 0, 0, 0, 0, 0, 0, -64, -64),
                (144, 14, 432, 400, -22, 0, 48, 0, 0, 0, 0, 0, 0, -64, -64),
                (144, 48, 432, -57, 80, 0, 48, 0, 0, 0, 0, 0, 0, -64, -64),
                (112, 16, 432, 304, -12, 80, 48, 0, 0, 0, 0, 0, 0, 0, 0),
                (144, 144, 432, 16, 144, 16, 48, 0, 0, 0, 0, 0, 0, 0, 0),
                (57, 36, -11, 368, 16, 68, 464, 0, 0, 0, 0, 0, 0, 0, 0),
                (144, 11, 176, -10, -45, 0, 16, 0, 0, 0, 0, 0, 0, -64, -64),
                (464, 14, 14, 57, -15, -54, 17, 0, 0, 0, 0, 0, 0, 0, 0),
                (48, 208, -12, 16, -57, 29, 80, 0, 0, 0, 0, 0, 0, 0, 0),
                (68, 272, 9, -65, -14, 272, 0, 0, 0, 0, 0, 0, 0, -64, -64),
                (144, -37, 176, -48, -14, 0, 16, 0, 0, 0, 0, 0, 0, -64, -64),
                (144, 33, -40, 336, 46, -55, -12, 0, 0, 0, 0, 0, 0, 0, 0),
                (80, 464, 16, 9, 14, 4, 208, 0, 0, 0, 0, 0, 0, 0, 0),
                (68, 272, 70, -65, -14, 0, -8, 0, 0, 0, 0, 0, 0, -64, -64),
                (-32, 16, -24, 13, -48, 176, 16, 0, 0, 0, 0, 0, 0, 0, 0),
                (144, 80, 176, 46, -5, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0),
                (464, 14, -18, -10, -10, 0, 432, 0, 0, 0, 0, 0, 0, -64, -64),
                (32, 20, 46, 208, 48, 42, 144, 0, 0, 0, 0, 0, 0, 0, 0),
                (176, -59, 16, -60, -37, 0, 0, 0, 0, 0, 0, -64, -64, -64, -64),
                (-20, 16, 464, 0, 400, 16, 55, 0, 0, 0, 0, 0, 0, -64, -64),
                (68, 38, 70, 432, 46, 16, 74, 0, 0, 0, 0, 0, 0, 0, 0),
                (80, -56, 48, 12, -37, 5, 80, 0, 0, 0, 0, 0, 0, 0, 0),
                (400, -20, 22, 0, -19, 208, 57, 0, 0, 0, 0, 0, 0, -64, -64),
                (48, 176, -69, -4, 48, -71, -17, 0, 0, 0, 0, 0, 0, 0, 0),
                (1, 1, 2, -1, 112, 368, 38, 0, 0, 0, 0, 0, 0, 0, 0),
                (56, 55, 5, 46, 1, 3, 368, 0, 0, 0, 0, 0, 0, 0, 0),
                (176, 80, 16, 208, 60, 0, 0, 0, 0, 0, 0, -64, -64, -64, -64),
                (68, 32, 272, 20, 16, 176, 9, 0, 0, 0, 0, 0, 0, 0, 0),
                (112, -17, -4, 16, 2, -4, -1, 0, 0, 0, 0, 0, 0, 0, 0),
                (20, -75, -22, 0, 208, 208, 432, 0, 0, 0, 0, 0, 0, -64, -64),
                (-50, -51, -37, 12, 0, 12, -36, 0, 0, 0, 0, 0, 0, -64, -64),
                (56, 55, 5, 46, 48, 3, 112, 0, 0, 0, 0, 0, 0, 0, 0),
                (176, 1, 16, 1, 2, 0, 0, 0, 0, 0, 0, -64, -64, -64, -64),
                (16, -42, 42, -70, -38, 144, 46, 0, 0, 0, 0, 0, 0, 0, 0),
                (-9, 176, -9, -13, -15, -9, 432, 0, 0, 0, 0, 0, 0, 0, 0),
                (21, 432, 208, 16, 7, 0, -22, 0, 0, 0, 0, 0, 0, -64, -64),
                (9, 9, 208, 8, -37, 112, 9, 0, 0, 0, 0, 0, 0, 0, 0),
                (80, 208, -5, -48, 0, 80, -4, 0, 0, 0, 0, 0, 0, -64, -64),
                (-32, 400, -24, -7, 144, 368, 400, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 2, 4, 7, -5, 0, 304, 0, 0, 0, 0, 0, 0, -64, -64),
                (112, 144, -4, 16, 432, -4, -4, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 17, 16, 13, 16, 34, 46, 0, 0, 0, 0, 0, 0, 0, 0),
                (-17, 16, -16, -19, 8, 0, -16, 0, 0, 0, 0, 0, 0, -64, -64),
                (464, -58, 11, 80, -57, -54, 13, 0, 0, 0, 0, 0, 0, 0, 0),
                (17, 17, 48, 48, 432, -48, 30, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, -7, 13, -8, -7, 48, 15, 0, 0, 0, 0, 0, 0, 0, 0),
                (176, 42, 16, 144, 46, 0, 0, 0, 0, 0, 0, -64, -64, -64, -64),
                (-32, -32, 400, 16, 0, 2, 4, 0, 0, 0, 0, 0, 0, -64, -64),
                (272, -17, -4, 80, -16, 16, 34, 0, 0, 0, 0, 0, 0, 0, 0),
                (-48, -8, -48, -8, -7, 0, -48, 0, 0, 0, 0, 0, 0, -64, -64)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((0, 0, 0, 0, 0, 0, 0, 18, 11, 12, -7, 2, -9, -6, -14),
                (0, 0, 0, 0, 0, 0, 0, 14, 9, 9, -2, -3, -11, -6, -12),
                (0, 0, 0, 0, 0, 0, 0, 12, 7, 8, -7, 4, -7, -4, -9),
                (0, 0, 0, 0, 0, 0, 0, 11, 6, -9, 7, 2, -6, -5, -11),
                (0, 0, 0, 0, 0, 0, 0, 10, -4, 8, -4, 6, -3, -3, -8),
                (0, 0, 0, 0, 0, 0, 0, 10, -1, 8, 1, 0, -5, 0, -6),
                (0, 0, 0, 0, 0, 0, 0, 9, -1, 6, -2, 1, -4, 0, -10),
                (0, 0, 0, 0, 0, 0, 0, 10, 1, 6, -4, 0, -6, 11, 5),
                (0, 0, 0, 0, 0, 0, 0, 8, 0, 3, -8, 4, -2, -1, -4),
                (0, 0, 0, 0, 0, 0, 0, 8, 1, 1, 10, 5, -2, -8, 10),
                (0, 0, 0, 0, 0, 10, 0, 6, -1, 1, -2, 5, -2, 10, 10),
                (0, 0, 0, 0, 0, 9, 0, 2, -1, -12, -5, 5, -2, 9, 9),
                (0, 0, 0, 0, 0, 9, 0, 8, 1, 0, -4, 4, -1, 9, 9),
                (0, 0, 0, 0, 0, 0, 0, 8, -2, -13, 2, 0, -8, -1, -7),
                (0, 0, 0, 0, 0, 0, 0, 3, 0, -1, -6, 5, 9, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, 2, -1, 3, -7, -8, 4, 9, -6),
                (0, 0, 0, 0, 0, 9, 0, -3, 1, -9, -2, -5, 6, 9, 9),
                (0, 0, 0, 0, 0, 0, 0, 1, 6, -9, -2, 3, -3, 17, -5),
                (0, 0, 0, 0, 0, 0, 0, 7, 1, 10, 0, -5, -11, 0, -8),
                (0, 0, 0, 0, 0, 0, -1, 8, 0, -8, -2, 5, 14, -1, -1),
                (0, 0, 0, 0, 0, 8, 0, 1, -7, 2, 0, -5, 5, 8, 8),
                (0, 0, 0, 0, 0, 0, 0, 3, 0, -7, 3, -1, -9, 2, -1),
                (0, 0, 0, 0, 0, 0, 0, 1, -2, -2, 4, 3, -6, -9, 3),
                (0, 0, 0, 0, 0, 10, 0, 6, 0, -7, -2, -3, 6, 10, 10),
                (0, 0, 0, 0, 0, 0, 0, 3, -8, 0, -6, 4, 16, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, -9, -2, 9, 4, -2, 6),
                (0, 0, 0, 0, 0, 10, 0, -2, 1, -6, 0, -1, -7, 10, 10),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, 7, 1, -1, -11, 3, -5),
                (0, 0, 0, 0, 0, -2, 8, 1, 12, -2, 0, -2, -2, 8, 8),
                (0, 0, 0, 8, 0, 0, 0, -11, -4, 1, 0, -1, -7, 8, 8),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, -5, 1, 3, 10, 0, 6),
                (0, 0, 0, 0, 0, 0, 0, 4, -6, -2, 0, -3, -15, 3, -4),
                (0, 0, 0, -10, 0, 0, 0, 10, 0, -10, -2, 6, -2, -10, -10),
                (0, 0, 0, 0, 0, 0, 0, 0, 4, 0, -7, 0, 10, -4, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 14, -14, -2, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, -5, -15, 3, -11, 9, -3),
                (0, 0, 0, 0, 0, -2, 8, 0, -9, -4, 4, -2, -2, 8, 8),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, 2, -2, 5, -5, 9, -1),
                (0, 0, 0, 0, 0, 0, 0, 4, -3, 6, 1, 0, 8, -2, 0),
                (0, 0, 0, 8, 0, 0, 0, 0, -1, -3, 8, -9, -3, 8, 8),
                (0, 0, 0, 0, 13, 0, 0, 2, -6, -3, 5, 10, 0, 13, 13),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, -11, 0, 2, -8, 8, -2),
                (0, 0, 0, 0, 0, -2, 8, 0, 5, -3, 0, -2, -2, 8, 8),
                (0, 0, 0, 0, 0, 0, 0, -7, 6, -10, 1, 0, 2, -7, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, -9, -2, 0, 16, 0, -1),
                (0, 0, 0, 0, 0, -9, 0, 0, 3, -3, 3, 5, -3, -9, -9),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, -7, 8, -1, -13, -11, 0),
                (0, 0, 0, 0, -7, 0, 0, 1, 0, 4, -10, 10, -2, -7, -7),
                (0, 0, 0, 0, 0, 0, 0, -6, -1, 3, -5, 7, 1, 1, -1),
                (0, 0, 0, 0, 0, 12, 0, 0, -2, 0, -9, -1, 1, 12, 12),
                (0, 0, 0, 0, 0, 0, 0, 5, 1, -3, 3, 0, 6, -10, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 6, 1, -9, 3, -4, 0),
                (0, 0, 0, 0, 0, 11, 0, 13, -1, -1, -8, -7, 0, 11, 11),
                (0, 0, 0, 0, 0, 0, 0, 4, -1, -11, 0, -7, -1, 7, -4),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 10, -2, 12, -1, -8, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 7, -14, -2, 0, 6, -4, 0),
                (0, 0, 0, 0, 0, -2, 7, 0, 2, -5, 0, -2, -2, 7, 7),
                (0, 0, 0, 0, -16, 0, 0, 2, -1, 3, 0, -2, 1, -16, -16),
                (0, 0, 0, 0, 0, 0, 0, 1, -9, 11, 0, 5, -1, -2, 4),
                (0, 0, 0, 0, 0, -12, 0, -2, -13, 18, 1, 9, 0, -12, -12)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;