LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE ieee.math_real.ALL;

LIBRARY work;
USE work.emp_data_types.ALL;
USE work.emp_device_decl.ALL;
USE work.kfout_data_formats.ALL;
USE work.kfout_config.ALL;

use work.hybrid_tools.all;
USE work.hybrid_config.ALL;
USE work.hybrid_data_types.ALL;
USE work.hybrid_data_formats.ALL;

PACKAGE kfout_luts IS

CONSTANT FloatV0Bins : REALS(0 TO 511 ) := (550763520.000000,
137690880.000000,
61195944.000000,
34422720.000000,
22030540.000000,
15298986.000000,
11240072.000000,
8605680.000000,
6799549.500000,
5507635.000000,
4551764.500000,
3824746.500000,
3258955.750000,
2810018.000000,
2447837.750000,
2151420.000000,
1905756.125000,
1699887.375000,
1525660.750000,
1376908.750000,
1248896.875000,
1137941.125000,
1041140.875000,
956186.625000,
881221.625000,
814738.937500,
755505.500000,
702504.500000,
654891.187500,
611959.437500,
573115.000000,
537855.000000,
505751.625000,
476439.031250,
449602.875000,
424971.843750,
402310.812500,
381415.187500,
362106.187500,
344227.187500,
327640.406250,
312224.218750,
297871.031250,
284485.281250,
271981.968750,
260285.218750,
249327.078125,
239046.656250,
229389.218750,
220305.406250,
211750.671875,
203684.734375,
196071.031250,
188876.375000,
182070.578125,
175626.125000,
169517.859375,
163722.796875,
158219.906250,
152989.859375,
148014.921875,
143278.750000,
138766.312500,
134463.750000,
130358.226562,
126437.906250,
122691.804688,
119109.757812,
115682.320312,
112400.718750,
109256.796875,
106242.960938,
103352.132812,
100577.703125,
97913.515625,
95353.796875,
92893.156250,
90526.546875,
88249.242188,
86056.796875,
83945.054688,
81910.101562,
79948.250000,
78056.054688,
76230.242188,
74467.757812,
72765.687500,
71121.320312,
69532.070312,
67995.492188,
66509.296875,
65071.304688,
63679.445312,
62331.769531,
61026.429688,
59761.664062,
58535.816406,
57347.304688,
56194.625000,
55076.351562,
53991.128906,
52937.667969,
51914.742188,
50921.183594,
49955.875000,
49017.757812,
48105.816406,
47219.093750,
46356.664062,
45517.644531,
44701.203125,
43906.531250,
43132.863281,
42379.464844,
41645.632812,
40930.699219,
40234.019531,
39554.976562,
38892.980469,
38247.464844,
37617.890625,
37003.730469,
36404.488281,
35819.687500,
35248.863281,
34691.578125,
34147.406250,
33615.937500,
33096.781250,
32589.556641,
32093.906250,
31609.476562,
31135.933594,
30672.951172,
30220.220703,
29777.439453,
29344.318359,
28920.580078,
28505.953125,
28100.179688,
27703.007812,
27314.199219,
26933.517578,
26560.740234,
26195.648438,
25838.033203,
25487.691406,
25144.425781,
24808.048828,
24478.378906,
24155.234375,
23838.449219,
23527.853516,
23223.289062,
22924.599609,
22631.636719,
22344.253906,
22062.310547,
21785.669922,
21514.199219,
21247.773438,
20986.263672,
20729.552734,
20477.525391,
20230.064453,
19987.062500,
19748.414062,
19514.013672,
19283.761719,
19057.560547,
18835.316406,
18616.939453,
18402.335938,
18191.421875,
17984.115234,
17780.330078,
17579.990234,
17383.017578,
17189.335938,
16998.873047,
16811.560547,
16627.324219,
16446.101562,
16267.826172,
16092.432617,
15919.861328,
15750.050781,
15582.942383,
15418.479492,
15256.607422,
15097.270508,
14940.416016,
14785.994141,
14633.954102,
14484.247070,
14336.826172,
14191.643555,
14048.656250,
13907.818359,
13769.087891,
13632.422852,
13497.782227,
13365.126953,
13234.416992,
13105.616211,
12978.685547,
12853.590820,
12730.295898,
12608.765625,
12488.968750,
12370.870117,
12254.439453,
12139.644531,
12026.454102,
11914.840820,
11804.773438,
11696.224609,
11589.166016,
11483.570312,
11379.411133,
11276.663086,
11175.300781,
11075.298828,
10976.632812,
10879.279297,
10783.215820,
10688.417969,
10594.866211,
10502.536133,
10411.408203,
10321.461914,
10232.674805,
10145.029297,
10058.504883,
9973.083008,
9888.744141,
9805.471680,
9723.245117,
9642.049805,
9561.866211,
9482.679688,
9404.472656,
9327.228516,
9250.932617,
9175.568359,
9101.122070,
9027.578125,
8954.921875,
8883.139648,
8812.215820,
8742.139648,
8672.894531,
8604.469727,
8536.851562,
8470.027344,
8403.984375,
8338.710938,
8274.195312,
8210.424805,
8147.389160,
8085.076660,
8023.476562,
7962.577148,
7902.369141,
7842.840820,
7783.983398,
7725.785156,
7668.237793,
7611.331055,
7555.055176,
7499.400879,
7444.359863,
7389.922363,
7336.079590,
7282.823242,
7230.145020,
7178.035645,
7126.488281,
7075.493652,
7025.044922,
6975.133301,
6925.751953,
6876.893555,
6828.549805,
6780.714355,
6733.379395,
6686.538574,
6640.185059,
6594.311523,
6548.912109,
6503.979980,
6459.508301,
6415.491211,
6371.922852,
6328.796387,
6286.106445,
6243.847168,
6202.012207,
6160.596680,
6119.594727,
6079.000488,
6038.808594,
5999.014160,
5959.612305,
5920.596680,
5881.963379,
5843.706543,
5805.822266,
5768.304688,
5731.149902,
5694.353027,
5657.909180,
5621.813965,
5586.063477,
5550.652832,
5515.577637,
5480.833984,
5446.417480,
5412.324219,
5378.549805,
5345.090820,
5311.943359,
5279.102539,
5246.565918,
5214.329102,
5182.388184,
5150.740234,
5119.381348,
5088.307617,
5057.516113,
5027.003418,
4996.765625,
4966.800293,
4937.103516,
4907.672363,
4878.503418,
4849.593750,
4820.940430,
4792.540039,
4764.390137,
4736.487793,
4708.829102,
4681.412598,
4654.234863,
4627.292480,
4600.583984,
4574.105957,
4547.855469,
4521.830566,
4496.028809,
4470.446777,
4445.082520,
4419.933594,
4394.997559,
4370.271973,
4345.754395,
4321.442383,
4297.333984,
4273.426758,
4249.718262,
4226.207031,
4202.890137,
4179.765625,
4156.831055,
4134.085449,
4111.525391,
4089.149902,
4066.956543,
4044.943115,
4023.108154,
4001.449463,
3979.965332,
3958.653564,
3937.512695,
3916.540527,
3895.735596,
3875.095947,
3854.619873,
3834.305664,
3814.151855,
3794.156250,
3774.317627,
3754.634033,
3735.104004,
3715.726074,
3696.498535,
3677.419922,
3658.488525,
3639.703125,
3621.061768,
3602.563477,
3584.206543,
3565.989502,
3547.910889,
3529.969727,
3512.164062,
3494.492676,
3476.954590,
3459.548096,
3442.271973,
3425.125000,
3408.105713,
3391.212891,
3374.445557,
3357.802246,
3341.281738,
3324.882812,
3308.604248,
3292.445068,
3276.404053,
3260.479736,
3244.671387,
3228.977783,
3213.397705,
3197.930176,
3182.573975,
3167.328125,
3152.191406,
3137.163330,
3122.242188,
3107.427246,
3092.717529,
3078.112061,
3063.609863,
3049.209717,
3034.911133,
3020.712646,
3006.613525,
2992.613037,
2978.710205,
2964.903809,
2951.193359,
2937.577637,
2924.056152,
2910.627686,
2897.291504,
2884.046631,
2870.892578,
2857.828125,
2844.852783,
2831.965576,
2819.165771,
2806.452637,
2793.825195,
2781.282715,
2768.824707,
2756.449951,
2744.158203,
2731.948242,
2719.819824,
2707.771973,
2695.803955,
2683.915039,
2672.104492,
2660.372070,
2648.716553,
2637.137451,
2625.634033,
2614.205811,
2602.852051,
2591.572266,
2580.365479,
2569.231201,
2558.168701,
2547.177734,
2536.257324,
2525.407227,
2514.626221,
2503.914307,
2493.270752,
2482.694824,
2472.186035,
2461.743896,
2451.367920,
2441.057129,
2430.811279,
2420.629883,
2410.512451,
2400.458008,
2390.466553,
2380.537354,
2370.669922,
2360.863525,
2351.118164,
2341.432617,
2331.807129,
2322.240723,
2312.733154,
2303.283691,
2293.892090,
2284.557861,
2275.280518,
2266.059570,
2256.894531,
2247.784912,
2238.730469,
2229.730469,
2220.784912,
2211.892822,
2203.053955,
2194.268311,
2185.534912,
2176.853516,
2168.223633,
2159.645264,
2151.117432,
2142.640137,
2134.212891,
2125.835205,
2117.506836,
2109.227295,
2100.996094  );

CONSTANT FloatV1Bins : REALS(0 TO 1023 ) := ( 625.663757,
156.415939,
69.518196,
39.103985,
25.026550,
17.379549,
12.768648,
9.775996,
7.724244,
6.256638,
5.170775,
4.344887,
3.702152,
3.192162,
2.780728,
2.443999,
2.164927,
1.931061,
1.733141,
1.564159,
1.418739,
1.292694,
1.182729,
1.086222,
1.001062,
0.925538,
0.858249,
0.798041,
0.743952,
0.695182,
0.651055,
0.611000,
0.574531,
0.541232,
0.510746,
0.482765,
0.457022,
0.433285,
0.411350,
0.391040,
0.372197,
0.354685,
0.338380,
0.323173,
0.308970,
0.295682,
0.283234,
0.271555,
0.260585,
0.250266,
0.240547,
0.231385,
0.222735,
0.214562,
0.206831,
0.199510,
0.192571,
0.185988,
0.179737,
0.173795,
0.168144,
0.162764,
0.157638,
0.152750,
0.148086,
0.143633,
0.139377,
0.135308,
0.131414,
0.127686,
0.124115,
0.120691,
0.117407,
0.114256,
0.111229,
0.108321,
0.105526,
0.102838,
0.100251,
0.097760,
0.095361,
0.093049,
0.090821,
0.088671,
0.086597,
0.084595,
0.082661,
0.080793,
0.078988,
0.077242,
0.075554,
0.073921,
0.072339,
0.070808,
0.069326,
0.067889,
0.066496,
0.065146,
0.063837,
0.062566,
0.061334,
0.060137,
0.058975,
0.057846,
0.056750,
0.055684,
0.054648,
0.053641,
0.052661,
0.051708,
0.050780,
0.049878,
0.048999,
0.048143,
0.047309,
0.046497,
0.045706,
0.044934,
0.044182,
0.043449,
0.042734,
0.042036,
0.041355,
0.040691,
0.040042,
0.039409,
0.038791,
0.038187,
0.037598,
0.037022,
0.036458,
0.035908,
0.035370,
0.034844,
0.034330,
0.033827,
0.033335,
0.032854,
0.032383,
0.031922,
0.031470,
0.031029,
0.030596,
0.030173,
0.029758,
0.029352,
0.028954,
0.028564,
0.028182,
0.027807,
0.027440,
0.027080,
0.026727,
0.026382,
0.026042,
0.025709,
0.025383,
0.025063,
0.024748,
0.024440,
0.024137,
0.023840,
0.023549,
0.023262,
0.022981,
0.022705,
0.022434,
0.022168,
0.021906,
0.021649,
0.021397,
0.021149,
0.020905,
0.020665,
0.020430,
0.020198,
0.019971,
0.019747,
0.019527,
0.019311,
0.019098,
0.018889,
0.018683,
0.018480,
0.018281,
0.018085,
0.017892,
0.017702,
0.017515,
0.017331,
0.017150,
0.016972,
0.016797,
0.016624,
0.016454,
0.016287,
0.016122,
0.015959,
0.015799,
0.015642,
0.015486,
0.015333,
0.015183,
0.015034,
0.014888,
0.014744,
0.014602,
0.014462,
0.014323,
0.014187,
0.014053,
0.013921,
0.013791,
0.013662,
0.013535,
0.013410,
0.013287,
0.013165,
0.013045,
0.012927,
0.012810,
0.012695,
0.012581,
0.012469,
0.012359,
0.012250,
0.012142,
0.012036,
0.011931,
0.011827,
0.011725,
0.011624,
0.011525,
0.011426,
0.011329,
0.011234,
0.011139,
0.011046,
0.010953,
0.010862,
0.010772,
0.010683,
0.010596,
0.010509,
0.010423,
0.010339,
0.010255,
0.010173,
0.010091,
0.010011,
0.009931,
0.009852,
0.009775,
0.009698,
0.009622,
0.009547,
0.009473,
0.009399,
0.009327,
0.009255,
0.009185,
0.009115,
0.009045,
0.008977,
0.008909,
0.008843,
0.008776,
0.008711,
0.008646,
0.008582,
0.008519,
0.008457,
0.008395,
0.008334,
0.008273,
0.008213,
0.008154,
0.008096,
0.008038,
0.007980,
0.007924,
0.007868,
0.007812,
0.007757,
0.007703,
0.007649,
0.007596,
0.007543,
0.007491,
0.007440,
0.007388,
0.007338,
0.007288,
0.007238,
0.007189,
0.007141,
0.007093,
0.007045,
0.006998,
0.006952,
0.006906,
0.006860,
0.006815,
0.006770,
0.006726,
0.006682,
0.006638,
0.006595,
0.006553,
0.006511,
0.006469,
0.006427,
0.006386,
0.006346,
0.006306,
0.006266,
0.006226,
0.006187,
0.006148,
0.006110,
0.006072,
0.006034,
0.005997,
0.005960,
0.005923,
0.005887,
0.005851,
0.005816,
0.005780,
0.005745,
0.005711,
0.005676,
0.005642,
0.005609,
0.005575,
0.005542,
0.005509,
0.005477,
0.005444,
0.005412,
0.005381,
0.005349,
0.005318,
0.005287,
0.005257,
0.005226,
0.005196,
0.005166,
0.005137,
0.005107,
0.005078,
0.005050,
0.005021,
0.004993,
0.004965,
0.004937,
0.004909,
0.004882,
0.004855,
0.004828,
0.004801,
0.004774,
0.004748,
0.004722,
0.004696,
0.004671,
0.004645,
0.004620,
0.004595,
0.004570,
0.004546,
0.004521,
0.004497,
0.004473,
0.004449,
0.004426,
0.004402,
0.004379,
0.004356,
0.004333,
0.004310,
0.004288,
0.004265,
0.004243,
0.004221,
0.004199,
0.004178,
0.004156,
0.004135,
0.004114,
0.004092,
0.004072,
0.004051,
0.004030,
0.004010,
0.003990,
0.003970,
0.003950,
0.003930,
0.003910,
0.003891,
0.003872,
0.003852,
0.003833,
0.003814,
0.003796,
0.003777,
0.003759,
0.003740,
0.003722,
0.003704,
0.003686,
0.003668,
0.003650,
0.003633,
0.003615,
0.003598,
0.003581,
0.003564,
0.003547,
0.003530,
0.003513,
0.003497,
0.003480,
0.003464,
0.003448,
0.003432,
0.003415,
0.003400,
0.003384,
0.003368,
0.003353,
0.003337,
0.003322,
0.003306,
0.003291,
0.003276,
0.003261,
0.003246,
0.003232,
0.003217,
0.003203,
0.003188,
0.003174,
0.003160,
0.003145,
0.003131,
0.003117,
0.003103,
0.003090,
0.003076,
0.003062,
0.003049,
0.003035,
0.003022,
0.003009,
0.002996,
0.002983,
0.002970,
0.002957,
0.002944,
0.002931,
0.002919,
0.002906,
0.002894,
0.002881,
0.002869,
0.002857,
0.002844,
0.002832,
0.002820,
0.002808,
0.002797,
0.002785,
0.002773,
0.002761,
0.002750,
0.002738,
0.002727,
0.002716,
0.002704,
0.002693,
0.002682,
0.002671,
0.002660,
0.002649,
0.002638,
0.002627,
0.002617,
0.002606,
0.002595,
0.002585,
0.002574,
0.002564,
0.002553,
0.002543,
0.002533,
0.002523,
0.002513,
0.002503,
0.002493,
0.002483,
0.002473,
0.002463,
0.002453,
0.002444,
0.002434,
0.002424,
0.002415,
0.002405,
0.002396,
0.002387,
0.002377,
0.002368,
0.002359,
0.002350,
0.002341,
0.002332,
0.002323,
0.002314,
0.002305,
0.002296,
0.002287,
0.002279,
0.002270,
0.002261,
0.002253,
0.002244,
0.002236,
0.002227,
0.002219,
0.002211,
0.002202,
0.002194,
0.002186,
0.002178,
0.002170,
0.002162,
0.002154,
0.002146,
0.002138,
0.002130,
0.002122,
0.002114,
0.002106,
0.002099,
0.002091,
0.002083,
0.002076,
0.002068,
0.002061,
0.002053,
0.002046,
0.002039,
0.002031,
0.002024,
0.002017,
0.002009,
0.002002,
0.001995,
0.001988,
0.001981,
0.001974,
0.001967,
0.001960,
0.001953,
0.001946,
0.001939,
0.001932,
0.001926,
0.001919,
0.001912,
0.001906,
0.001899,
0.001892,
0.001886,
0.001879,
0.001873,
0.001866,
0.001860,
0.001853,
0.001847,
0.001841,
0.001834,
0.001828,
0.001822,
0.001816,
0.001810,
0.001803,
0.001797,
0.001791,
0.001785,
0.001779,
0.001773,
0.001767,
0.001761,
0.001755,
0.001750,
0.001744,
0.001738,
0.001732,
0.001726,
0.001721,
0.001715,
0.001709,
0.001704,
0.001698,
0.001693,
0.001687,
0.001681,
0.001676,
0.001670,
0.001665,
0.001660,
0.001654,
0.001649,
0.001644,
0.001638,
0.001633,
0.001628,
0.001622,
0.001617,
0.001612,
0.001607,
0.001602,
0.001597,
0.001591,
0.001586,
0.001581,
0.001576,
0.001571,
0.001566,
0.001561,
0.001557,
0.001552,
0.001547,
0.001542,
0.001537,
0.001532,
0.001527,
0.001523,
0.001518,
0.001513,
0.001509,
0.001504,
0.001499,
0.001495,
0.001490,
0.001485,
0.001481,
0.001476,
0.001472,
0.001467,
0.001463,
0.001458,
0.001454,
0.001449,
0.001445,
0.001441,
0.001436,
0.001432,
0.001428,
0.001423,
0.001419,
0.001415,
0.001411,
0.001406,
0.001402,
0.001398,
0.001394,
0.001390,
0.001385,
0.001381,
0.001377,
0.001373,
0.001369,
0.001365,
0.001361,
0.001357,
0.001353,
0.001349,
0.001345,
0.001341,
0.001337,
0.001333,
0.001330,
0.001326,
0.001322,
0.001318,
0.001314,
0.001310,
0.001307,
0.001303,
0.001299,
0.001295,
0.001292,
0.001288,
0.001284,
0.001281,
0.001277,
0.001273,
0.001270,
0.001266,
0.001262,
0.001259,
0.001255,
0.001252,
0.001248,
0.001245,
0.001241,
0.001238,
0.001234,
0.001231,
0.001227,
0.001224,
0.001220,
0.001217,
0.001214,
0.001210,
0.001207,
0.001204,
0.001200,
0.001197,
0.001194,
0.001190,
0.001187,
0.001184,
0.001181,
0.001177,
0.001174,
0.001171,
0.001168,
0.001164,
0.001161,
0.001158,
0.001155,
0.001152,
0.001149,
0.001146,
0.001143,
0.001139,
0.001136,
0.001133,
0.001130,
0.001127,
0.001124,
0.001121,
0.001118,
0.001115,
0.001112,
0.001109,
0.001106,
0.001103,
0.001101,
0.001098,
0.001095,
0.001092,
0.001089,
0.001086,
0.001083,
0.001080,
0.001078,
0.001075,
0.001072,
0.001069,
0.001066,
0.001064,
0.001061,
0.001058,
0.001055,
0.001053,
0.001050,
0.001047,
0.001044,
0.001042,
0.001039,
0.001036,
0.001034,
0.001031,
0.001028,
0.001026,
0.001023,
0.001021,
0.001018,
0.001015,
0.001013,
0.001010,
0.001008,
0.001005,
0.001003,
0.001000,
0.000997,
0.000995,
0.000992,
0.000990,
0.000987,
0.000985,
0.000983,
0.000980,
0.000978,
0.000975,
0.000973,
0.000970,
0.000968,
0.000965,
0.000963,
0.000961,
0.000958,
0.000956,
0.000954,
0.000951,
0.000949,
0.000947,
0.000944,
0.000942,
0.000940,
0.000937,
0.000935,
0.000933,
0.000930,
0.000928,
0.000926,
0.000924,
0.000921,
0.000919,
0.000917,
0.000915,
0.000913,
0.000910,
0.000908,
0.000906,
0.000904,
0.000902,
0.000900,
0.000897,
0.000895,
0.000893,
0.000891,
0.000889,
0.000887,
0.000885,
0.000883,
0.000880,
0.000878,
0.000876,
0.000874,
0.000872,
0.000870,
0.000868,
0.000866,
0.000864,
0.000862,
0.000860,
0.000858,
0.000856,
0.000854,
0.000852,
0.000850,
0.000848,
0.000846,
0.000844,
0.000842,
0.000840,
0.000838,
0.000836,
0.000834,
0.000832,
0.000830,
0.000829,
0.000827,
0.000825,
0.000823,
0.000821,
0.000819,
0.000817,
0.000815,
0.000813,
0.000812,
0.000810,
0.000808,
0.000806,
0.000804,
0.000802,
0.000801,
0.000799,
0.000797,
0.000795,
0.000793,
0.000792,
0.000790,
0.000788,
0.000786,
0.000785,
0.000783,
0.000781,
0.000779,
0.000778,
0.000776,
0.000774,
0.000772,
0.000771,
0.000769,
0.000767,
0.000766,
0.000764,
0.000762,
0.000761,
0.000759,
0.000757,
0.000756,
0.000754,
0.000752,
0.000751,
0.000749,
0.000747,
0.000746,
0.000744,
0.000742,
0.000741,
0.000739,
0.000738,
0.000736,
0.000734,
0.000733,
0.000731,
0.000730,
0.000728,
0.000727,
0.000725,
0.000723,
0.000722,
0.000720,
0.000719,
0.000717,
0.000716,
0.000714,
0.000713,
0.000711,
0.000710,
0.000708,
0.000707,
0.000705,
0.000704,
0.000702,
0.000701,
0.000699,
0.000698,
0.000696,
0.000695,
0.000693,
0.000692,
0.000690,
0.000689,
0.000687,
0.000686,
0.000685,
0.000683,
0.000682,
0.000680,
0.000679,
0.000677,
0.000676,
0.000675,
0.000673,
0.000672,
0.000670,
0.000669,
0.000668,
0.000666,
0.000665,
0.000664,
0.000662,
0.000661,
0.000660,
0.000658,
0.000657,
0.000655,
0.000654,
0.000653,
0.000651,
0.000650,
0.000649,
0.000647,
0.000646,
0.000645,
0.000644,
0.000642,
0.000641,
0.000640,
0.000638,
0.000637,
0.000636,
0.000635,
0.000633,
0.000632,
0.000631,
0.000629,
0.000628,
0.000627,
0.000626,
0.000624,
0.000623,
0.000622,
0.000621,
0.000619,
0.000618,
0.000617,
0.000616,
0.000615,
0.000613,
0.000612,
0.000611,
0.000610,
0.000609,
0.000607,
0.000606,
0.000605,
0.000604,
0.000603,
0.000601,
0.000600,
0.000599,
0.000598,
0.000597 );

--CONSTANT rescaledChi2RphiBins : REALS( 0 TO ( 2**widthChi2RPhi ) - 1 ) := ( 0.0, 206536098.38900286, 309804147.5835043, 413072196.7780057, 516340245.97250724, 619608295.1670086, 722876344.36151, 826144393.5560114, 1032680491.9450145, 1239216590.3340173, 2065360983.890029, 3098041475.835043, 4130721967.780058, 7228763443.615101, 12392165903.340172, 41307219677.800575);
CONSTANT rescaledChi2RphiBins : REALS( 0 TO (2**widthChi2RPhi) - 1 ) := ( 0.0, 22948455.376555875, 34422683.06483381, 45896910.75311175, 57371138.44138969, 68845366.12966762, 80319593.81794555, 91793821.5062235, 114742276.88277937, 137690732.25933525, 229484553.76555875, 344226830.64833814, 458969107.5311175, 803195938.1794556, 1376907322.5933526, 4589691075.311175 );
CONSTANT rescaledChi2RZBins : REALS( 0 TO ( 2**widthChi2RZ ) - 1 ) := (   0.0, 6308223.406369258, 12616446.812738515, 18924670.219107773, 25232893.62547703, 31541117.031846285, 37849340.43821555, 44157563.84458481, 50465787.25095406, 56774010.657323316, 63082234.06369257, 75698680.8764311, 100931574.50190812, 126164468.12738514, 252328936.25477028, 630822340.6369258);

END kfout_luts;