library ieee;
use ieee.std_logic_1164.all;



package tracklet_components is


component IR_PS10G_1_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS10G_2_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS10G_2_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS10G_3_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS10G_3_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS_1_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS_1_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS_2_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_PS_2_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_1_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0);
    hOutputStubs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_1_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_2_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_2_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_3_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_3_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_4_A
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component IR_2S_4_B
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    hInputStubs_V_dout : IN STD_LOGIC_VECTOR (38 downto 0);
    hInputStubs_V_empty_n : IN STD_LOGIC;
    hInputStubs_V_read : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    hLinkWord_V : IN STD_LOGIC_VECTOR (19 downto 0);
    hPhBnWord_V : IN STD_LOGIC_VECTOR (31 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    hOutputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    hOutputStubs_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0) );
end component;

component VMR_L1PHID
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    memoriesAS_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesAS_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0);
    memoriesTEI_0_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_0_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_0_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_0_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_0_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_0_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_0_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_0_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_0_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_0_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_0_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_0_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_0_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_0_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_0_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_0_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_1_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_1_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_1_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_1_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_1_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_1_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_1_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_1_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_1_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_1_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_1_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_1_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_1_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_1_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_1_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_1_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_2_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_2_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_2_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_2_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_2_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_2_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_2_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_2_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_2_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_2_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_2_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_2_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_2_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_2_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_2_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_2_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_3_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_3_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_3_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_3_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_3_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_3_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_3_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_3_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_3_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_3_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_3_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_3_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0);
    memoriesTEI_3_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEI_3_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEI_3_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEI_3_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (21 downto 0) );
end component;

component VMR_L2PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    memoriesAS_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesAS_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0);
    memoriesTEO_0_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_0_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_0_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_0_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_0_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_0_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_0_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_0_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_0_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_0_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_0_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_0_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_1_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_1_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_1_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_1_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_1_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_1_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_1_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_1_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_1_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_1_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_1_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_1_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_2_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_2_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_2_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_2_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_2_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_2_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_2_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_2_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_2_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_2_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_2_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_2_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_3_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_3_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_3_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_3_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_3_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_3_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_3_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_3_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_3_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_3_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_3_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_3_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_4_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_4_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_4_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_4_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_4_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_4_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_4_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_4_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_4_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_4_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_4_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_4_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_5_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_5_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_5_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_5_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_5_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_5_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_5_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_5_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_5_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_5_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_5_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_5_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_6_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_6_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_6_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_6_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_6_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_6_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_6_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_6_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_6_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_6_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_6_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_6_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_7_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_7_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_7_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_7_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_7_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_7_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_7_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_7_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesTEO_7_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    memoriesTEO_7_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesTEO_7_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesTEO_7_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0) );
end component;

component VMR_L3PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    memoriesAS_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesAS_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0);
    memoriesME_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesME_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesME_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesME_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesME_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesME_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesME_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0);
    memoriesME_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (15 downto 0) );
end component;

component VMR_L4PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    memoriesAS_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesAS_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0);
    memoriesME_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0) );
end component;

component VMR_L5PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    memoriesAS_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesAS_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0);
    memoriesME_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0) );
end component;

component VMR_L6PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputStubs_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubs_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    inputStubs_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputStubs_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    memoriesAS_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesAS_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesAS_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (35 downto 0);
    memoriesME_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0);
    memoriesME_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    memoriesME_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    memoriesME_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (16 downto 0) );
end component;

component TE_L1L2
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    instubinnerdata_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    instubinnerdata_dataarray_data_V_ce0 : OUT STD_LOGIC;
    instubinnerdata_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (21 downto 0);
    instubinnerdata_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    instubinnerdata_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    instubouterdata_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    instubouterdata_dataarray_data_V_ce0 : OUT STD_LOGIC;
    instubouterdata_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (15 downto 0);
    instubouterdata_nentries_0_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_0_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_0_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_0_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_0_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_0_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_0_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_0_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    instubouterdata_nentries_1_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    bendinnertable_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    bendinnertable_V_ce0 : OUT STD_LOGIC;
    bendinnertable_V_q0 : IN STD_LOGIC_VECTOR (0 downto 0);
    bendoutertable_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    bendoutertable_V_ce0 : OUT STD_LOGIC;
    bendoutertable_V_q0 : IN STD_LOGIC_VECTOR (0 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    outstubpair_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    outstubpair_dataarray_data_V_ce0 : OUT STD_LOGIC;
    outstubpair_dataarray_data_V_we0 : OUT STD_LOGIC;
    outstubpair_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (13 downto 0) );
end component;

component TC_L1L2F
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    innerStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    innerStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    innerStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    outerStubs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    outerStubs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    outerStubs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    stubPairs_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_4_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_5_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_6_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_7_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_8_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    stubPairs_8_dataarray_data_V_ce0 : OUT STD_LOGIC;
    stubPairs_8_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    stubPairs_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_4_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_4_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_5_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_5_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_6_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_6_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_7_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_7_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_8_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    stubPairs_8_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    trackletParameters_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    trackletParameters_dataarray_data_V_ce0 : OUT STD_LOGIC;
    trackletParameters_dataarray_data_V_we0 : OUT STD_LOGIC;
    trackletParameters_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (69 downto 0);
    projout_barrel_ps_13_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projout_barrel_ps_13_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projout_barrel_ps_13_dataarray_data_V_we0 : OUT STD_LOGIC;
    projout_barrel_ps_13_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (59 downto 0);
    projout_barrel_2s_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projout_barrel_2s_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projout_barrel_2s_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    projout_barrel_2s_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (57 downto 0);
    projout_barrel_2s_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projout_barrel_2s_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projout_barrel_2s_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    projout_barrel_2s_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (57 downto 0);
    projout_barrel_2s_9_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projout_barrel_2s_9_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projout_barrel_2s_9_dataarray_data_V_we0 : OUT STD_LOGIC;
    projout_barrel_2s_9_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (57 downto 0) );
end component;

component PR_L3PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    projin_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projin_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projin_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (59 downto 0);
    projin_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    projin_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    allprojout_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allprojout_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_we0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (59 downto 0);
    vmprojout_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0) );
end component;

component PR_L4PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    projin_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projin_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projin_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (57 downto 0);
    projin_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    projin_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    allprojout_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allprojout_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_we0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (57 downto 0);
    vmprojout_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0) );
end component;

component PR_L5PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    projin_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projin_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projin_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (57 downto 0);
    projin_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    projin_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    allprojout_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allprojout_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_we0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (57 downto 0);
    vmprojout_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0) );
end component;

component PR_L6PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    projin_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    projin_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    projin_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (57 downto 0);
    projin_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    projin_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    allprojout_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allprojout_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_we0 : OUT STD_LOGIC;
    allprojout_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (57 downto 0);
    vmprojout_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_1_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_2_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_3_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_4_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_5_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_6_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0);
    vmprojout_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    vmprojout_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_we0 : OUT STD_LOGIC;
    vmprojout_7_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (23 downto 0) );
end component;

component ME_L3PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    inputStubData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (15 downto 0);
    inputStubData_nentries_0_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputProjectionData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputProjectionData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputProjectionData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (23 downto 0);
    inputProjectionData_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputProjectionData_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    outputCandidateMatch_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    outputCandidateMatch_dataarray_data_V_ce0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_we0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (13 downto 0) );
end component;

component ME_L4PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    inputStubData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (16 downto 0);
    inputStubData_nentries_0_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputProjectionData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputProjectionData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputProjectionData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (23 downto 0);
    inputProjectionData_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputProjectionData_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    outputCandidateMatch_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    outputCandidateMatch_dataarray_data_V_ce0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_we0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (13 downto 0) );
end component;

component ME_L5PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    inputStubData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (16 downto 0);
    inputStubData_nentries_0_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputProjectionData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputProjectionData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputProjectionData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (23 downto 0);
    inputProjectionData_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputProjectionData_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    outputCandidateMatch_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    outputCandidateMatch_dataarray_data_V_ce0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_we0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (13 downto 0) );
end component;

component ME_L6PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    inputStubData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputStubData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (16 downto 0);
    inputStubData_nentries_0_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_0_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_1_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_2_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_3_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_4_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_5_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_6_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_0 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_1 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_2 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_3 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_4 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_5 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_6 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputStubData_nentries_7_V_7 : IN STD_LOGIC_VECTOR (4 downto 0);
    inputProjectionData_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    inputProjectionData_dataarray_data_V_ce0 : OUT STD_LOGIC;
    inputProjectionData_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (23 downto 0);
    inputProjectionData_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    inputProjectionData_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    outputCandidateMatch_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    outputCandidateMatch_dataarray_data_V_ce0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_we0 : OUT STD_LOGIC;
    outputCandidateMatch_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (13 downto 0) );
end component;

component MC_L3PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    match_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_4_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_5_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_6_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_7_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    allstub_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allstub_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allstub_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    allproj_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allproj_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allproj_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (59 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    fullmatch_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (51 downto 0) );
end component;

component MC_L4PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    match_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_4_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_5_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_6_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_7_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    allstub_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allstub_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allstub_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    allproj_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allproj_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allproj_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (57 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    fullmatch_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (51 downto 0) );
end component;

component MC_L5PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    match_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_4_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_5_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_6_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_7_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    allstub_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allstub_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allstub_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    allproj_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allproj_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allproj_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (57 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    fullmatch_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (51 downto 0) );
end component;

component MC_L6PHIB
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    match_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_4_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_4_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_4_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_5_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_5_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_5_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_6_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_6_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_6_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_7_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    match_7_dataarray_data_V_ce0 : OUT STD_LOGIC;
    match_7_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (13 downto 0);
    match_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_4_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_5_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_6_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    match_7_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    allstub_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allstub_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allstub_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (35 downto 0);
    allproj_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    allproj_dataarray_data_V_ce0 : OUT STD_LOGIC;
    allproj_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (57 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    fullmatch_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_we0 : OUT STD_LOGIC;
    fullmatch_0_dataarray_data_V_d0 : OUT STD_LOGIC_VECTOR (51 downto 0) );
end component;

component FT_L1L2
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    bx_V : IN STD_LOGIC_VECTOR (2 downto 0);
    trackletParameters_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (9 downto 0);
    trackletParameters_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    trackletParameters_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (69 downto 0);
    barrelFullMatches_0_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    barrelFullMatches_0_dataarray_data_V_ce0 : OUT STD_LOGIC;
    barrelFullMatches_0_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (51 downto 0);
    barrelFullMatches_1_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    barrelFullMatches_1_dataarray_data_V_ce0 : OUT STD_LOGIC;
    barrelFullMatches_1_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (51 downto 0);
    barrelFullMatches_2_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    barrelFullMatches_2_dataarray_data_V_ce0 : OUT STD_LOGIC;
    barrelFullMatches_2_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (51 downto 0);
    barrelFullMatches_3_dataarray_data_V_address0 : OUT STD_LOGIC_VECTOR (7 downto 0);
    barrelFullMatches_3_dataarray_data_V_ce0 : OUT STD_LOGIC;
    barrelFullMatches_3_dataarray_data_V_q0 : IN STD_LOGIC_VECTOR (51 downto 0);
    barrelFullMatches_0_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    barrelFullMatches_0_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    barrelFullMatches_1_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    barrelFullMatches_1_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    barrelFullMatches_2_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    barrelFullMatches_2_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    barrelFullMatches_3_nentries_0_V : IN STD_LOGIC_VECTOR (6 downto 0);
    barrelFullMatches_3_nentries_1_V : IN STD_LOGIC_VECTOR (6 downto 0);
    bx_o_V : OUT STD_LOGIC_VECTOR (2 downto 0);
    bx_o_V_ap_vld : OUT STD_LOGIC;
    trackWord_V_din : OUT STD_LOGIC_VECTOR (83 downto 0);
    trackWord_V_full_n : IN STD_LOGIC;
    trackWord_V_write : OUT STD_LOGIC;
    barrelStubWords_0_V_din : OUT STD_LOGIC_VECTOR (45 downto 0);
    barrelStubWords_0_V_full_n : IN STD_LOGIC;
    barrelStubWords_0_V_write : OUT STD_LOGIC;
    barrelStubWords_1_V_din : OUT STD_LOGIC_VECTOR (45 downto 0);
    barrelStubWords_1_V_full_n : IN STD_LOGIC;
    barrelStubWords_1_V_write : OUT STD_LOGIC;
    barrelStubWords_2_V_din : OUT STD_LOGIC_VECTOR (45 downto 0);
    barrelStubWords_2_V_full_n : IN STD_LOGIC;
    barrelStubWords_2_V_write : OUT STD_LOGIC;
    barrelStubWords_3_V_din : OUT STD_LOGIC_VECTOR (45 downto 0);
    barrelStubWords_3_V_full_n : IN STD_LOGIC;
    barrelStubWords_3_V_write : OUT STD_LOGIC );
end component;


end;